TranslationLanguage=Svenska

"Remote to local path mappings.~Examples:~/share=\\pch\share~/var/downloads/music=Z:\music"="Mappning fjärr- till lokala sökvägar.~Till exempel:~/share=\\pch\share~/var/downloads/musik=Z:\musik"
%d x %s (have %d)=%d x %s (har %d)
%ds=%ds
%s (%d hashfails)=%s (%d hashfel)
%s (%s done)=%s (%s klar)
'%s' has finished downloading='%s' är klar med nedladdningen
%s%s%d downloading, %d seeding%s%s, %s=%s%s%d laddar ner, %d delar%s%s, %s
&All=&Alla
&Close=&Stäng
&Help=&Hjälp
&Ignore=&Ignorera
&No=&Nej
&OK=&OK
&Open=&Öppna
&Retry=&Försök igen
&Save=&Spara
&Unlock=Lås upp
&Yes=&Ja
/s=/s
Abort=Avbryt
About=Om
Active=Aktiv
Add new torrent=Lägg till ny torrent
&Add torrent=Lägg till torrent
Added on=Lades till
Are you sure to remove torrent '%s' and all associated DATA?=Är du säker på att du vill ta bort '%s' och all tillhörande data?
Are you sure to remove torrent '%s'?=Är du säker på att du vill ta bort torrenten '%s'?
Authentication=Autentisering
b=b
Cancel=Avbryt
Client=Klient
Close to tray=Stäng till aktivitetsfältet
Comment=Kommentar
Completed on=Avslutad den
Completed=Avslutad
Confirmation=Bekräftelse
connected=ansluten
Connecting to daemon=Ansluter till server
Connection error occurred=Anslutningsfel har inträffat
Copy=Kopiera
Country=Land
Created on=Skapad
D: %s/s=D: %s/s
Destination folder=Destinationsmapp
Disconnected=Frånkopplad
Donate to support further development=Donera för att stödja fortsatt utveckling
Donate via PayPal,WebMoney,Credit card=Donera via PayPal,WebMoney,Credit card
Done=Färdig
Don't download=Ladda inte ner
Down limit=Nedladdningsgräns
Down speed=Nedladdningshastighet
Down=Ner
Download complete=Nedladdning klar
Download speed=Nedladdingshastighet
Downloaded=Nedladdad
Downloading=Laddar ner
Enable DHT=Aktivera DHT
Enable Peer Exchange=Aktivera Peer Exchange
Enable port forwarding=Aktivera portvidarebefordran
Encryption disabled=Kryptering avstängt
Encryption enabled=Kryptering aktiverat
Encryption required=Kryptering krävs
Encryption=Kryptering
Error=Fel
ETA=ETA
E&xit=Avsluta
File name=Filnamn
Files=Filer
Finished=Färdig
Flag images archive is needed to display country flags.~Download this archive now?=Ett arkiv med flaggbilder är nödvändigt för att visa landsflaggor.~Vill du ladda ner denna nu?
Flags=Flaggor
GB=GB
General=Allmänt
Geo IP database is needed to resolve country by IP address.~Download this database now?=En geo-IP databas är nödvändig för att visa vilket land en IP-adress tillhör.~Önskar du att ladda ner denna databasen nu??
Global bandwidth settings=Global bredbands inställningar
Global peer limit=Max antal globala kamrater
Hash=Hash
Have=Har
Hide=Dölj
High priority=Hög prioritet
high=hög
Host=Värd
in swarm=i svärm
Inactive=Inaktiv
Incoming port is closed. Check your firewall settings=Inkommande port är stängd. Kontrollera brandväggs inställningarna
Incoming port tested successfully=Inkommande port är öppen
Incoming port=Inkommande port
Information=Information
KB/s=KB/s
KB=KB
Language=Språk
Last active=Senast aktiv
License=Licens
Low priority=Låg prioritet
low=låg
Max peers=Max antal peers
Maximum download speed=Max nedladdningshastighet
Maximum upload speed=Max uppladdningshastighet
MB=MB
Minimize to tray=Minimera till aktivitetsfältet
Name=Namn
No host name specified=Inget värdnamn specifierat
No proxy server specified=Ingen proxyserver specifierad
No to all=Nej till alla
Normal priority=Normal prioritet
normal=normal
of=av
Open containing folder=Öppna målmapp
Open=Öppna
Password=Lösenord
Paths=Sökvägar
Peer limit=Peer begränsning
Peers=Peers
Pieces=Delar
Port=Port
Priority=Prioritet
Properties=Egenskaper
Proxy password=Proxylösenord
Proxy port=Proxyport
Proxy server=Proxyserver
Proxy user name=Proxyanvändarnamn
Ratio=Förhållande
Reconnect in %d seconds=Anslut på nytt om %d sekunder
Remaining=Återstående
Remote host=Fjärrserver
Remove torrent and Data=Ta bort torrent och data
Remove torrent=Ta bort torrent
Remove=Ta bort
Resolve country=Check land
Resolve host name=Check värdnamn
seconds=sekunder
Seed ratio=Delningsförhållande
Seeding=Delar
Seeds=Delare
Select a .torrent to open=Välj en .torrent att öppna
Select all=Välj alla
Select none=Välj ingen
Setup columns=Ställ in kolumner
Share ratio=Delningsförhållande
Show country flag=Visa flagga
Show=Visa
Size=Storlek
skip=hoppa över
Start all torrents=Starta alla torrents
Start torrent=Starta torrent
Start=Starta
Status=Status
Stop all torrents=Stoppa alla torrents
Stop all=Stoppa alla
Stop torrent=Stoppa torrent
Stop=Stoppa
Stopped=Stoppad
TB=TB
Test port=Testa porten
T&ools=Verktyg
Torrent contents=Innehåll i torrent
Torrent properties=Egenskaper för torrent
Torrent verification may take a long time.~Are you sure to start verification of torrent '%s'?=Torrentverifikation kan ta lång tid.~Är du säker på att du vill starta torrentverifikation '%s'?
&Torrent=Torrent
Torrents (*.torrent)|*.torrent|All files (*.*)|*.*=Torrenter (*.torrent)|*.torrent|Alla filar (*.*)|*.*
Total size=Total storlek
Tracker status=Trackerstatus
Tracker update on=Tracker uppdaterad den
Tracker=Tracker
Trackers=Trackers
Transfer=Överföring
Transmission options=Alternativ för Transmission
Transmission%s at %s:%s=Transmission%s på %s:%s
Tray icon always visible=Ikon i aktivitetsfältet alltid synlig
Tray icon=Ikon i aktivitetsfältet
U: %s/s=U: %s/s
Unable to extract flag image=Kunde inte hämta flaggbild
Unable to get files list=Kunde inte hämta fillista
Unknown=Okänt
Up limit=Uppladdningsgräns
Up speed=Uppladdningshastighet
Up=Upp
Update complete=Uppdatering genomförd
Update GeoIP database=Uppdatera GeoIP-databas
Update in=Uppdaterar om
Updating=Uppdaterar
Upload speed=Uppladdningshastighet
Uploaded=Uppladdat
User name=Användarnamn
Verify torrent=Verifiera torrents
&Verify=Verifiera
Verifying=Verifierar
Version %s=Version %s
Waiting=Väntar
Warning=Varning
Wasted=Bortkastat
Working=Arbetar
Yes to &All=Ja till &allt
No tracker=Ingen tracker
%s downloaded=%s nedladdat
%s of %s downloaded=%s av %s nedladdat
%d torrents=%d torrents
Add .part extension to incomplete files=Lägg till .part på ofullständiga filer
Add torrent link=Lägg till en torrentlänk
Are you sure to remove %d selected torrents and all their associated DATA?=är du säker på att du önskar att ta bort %d valda torrenter och alla tilhörande data?
Are you sure to remove %d selected torrents?=är du säker på att du önskar att ta bort %d valda torrenter?
Bandwidth=Bandbredd
Directory for incomplete files=Mapp för ofullständiga filer
Download=Ladda ner
Enable blocklist=Aktivera blockeringslistan
ID=ID
Move torrent data from current location to new location=Flytta data från nuvarande plats till en ny plats
New location for torrent data=Ny plats för torrent data
No link was specified=Ingen länk specifierad
No torrent location was specified=Ingen torrentplats var specifierad
Path=Sökväg
Reannounce (get more peers)=Tillkännage (skaffa flera peers)
Set data location=Sätt dataplats
Size to download=Storlek på nedladdning
The block list has been updated successfully.~The list entries count: %d=Blockeringslistan blev uppdaterad.~Det är %d registrerade i listan
The directory for incomplete files was not specified=Mappen för ofullständiga filer var inte specifierad
The downloads directory was not specified=Nedladdningsmappen var inte specificerad
Torrent data location=Dataplats for torrent
Torrents=Torrents
Unable to execute "%s"=Kunde inte köra "%s"
Update blocklist=Uppdatera blockeringslista
URL of a .torrent file or a magnet link=Adressen till en .torrent-fil eller en magnet-länk
Columns setup=Kolumninställning
Add torrent=Lägg till torrent
Delete a .torrent file after a successful addition=Ta bort .torrent-filen efter den lagts till
Torrent=Torrent
Torrents verification may take a long time.~Are you sure to start verification of %d torrents?=Dataverifiering kan ta lång tid.~Är du säker på att du önskar att verifiera %d torrenter?
Unable to load OpenSSL library files: %s and %s=Klarade inte att ladda OpenSSL biblioteks filerna: %s och %s från OpenSSL
Use SSL=Använd SSL
Add tracker=Lägg till tracker
Alternate bandwidth settings=Alternativa bandbreddsinställingar
Apply alternate bandwidth settings automatically=Använd alternativa bandbreddsinställningar automatiskt
Are you sure to delete connection '%s'?=Är du säker på att du vill ta bort anslutningen '%s'?
Are you sure to remove tracker '%s'?=Är du säker på att du vill ta bort trackern '%s'?
Days=Dagar
Delete=Ta bort
Disk cache size=Storlek på diskcachen
  Download speeds (KB/s)=Nedladdingshastighet (KB/s)
Edit tracker=Redigera tracker
Enable Local Peer Discovery=Aktivera Lokal Peer-upptäckt
Free disk space=Ledigt diskutrymme
Free: %s=Ledigt: %s
From=Från
minutes=minuter
Misc=Diverse
New connection=Ny anslutning
New=Ny
No tracker URL was specified=Ingen trackeradress var specifierad
Proxy=Proxy
Remove tracker=Ta bort tracker
Rename=Byt namn
Speed limit menu items=Hastighetsbegränsningar
Stop seeding when inactive for=Avsluta delning när inaktiv i
The invalid time value was entered=Ett ogiltig tidsvärde angavs
to=till
Tracker announce URL=Trackerns annonseringsadress
Tracker properties=Trackerinställningar
Unlimited=Obegränsat
Upload speeds (KB/s)=Uppladdningshastighet (KB/s)
Use alternate bandwidth settings=Använd alternativa bandbreddsinställningar
average=genomsnitt
Browse=Bläddra
Enable µTP=Aktivera µTP
Select a folder for download=Välj nedladdningsmapp
Select torrent location=Välj torrentplats
A new version of %s is available.~Your current version: %s~The new version: %s~Do you wish to open the Downloads web page?=A new version of %s is available.~Your current version: %s~The new version: %s~Do you wish to open the Downloads web page?
Advanced=Avancerad
Check for new version every=Sök efter nya versioner varje
Check for updates=Sök efter uppdateringar
Consider active torrents as stalled when idle for=Anse att aktiva torrents är inaktiva efter
Do you wish to enable automatic checking for a new version of %s?=Vill du aktivera automatisk kontroll av nya versioner av %s?
Donate!=Donera!
Download queue size=Storlek på nedladdningskön
Error checking for new version=Fel vid koll efter ny version
Folder grouping=Gruppering av mappar
Force start=Tvångsstarta
Home page=Hemsida
Modify trackers=Ändra trackers
Move bottom=Flytta till botten av kön
Move down queue=Flytta ner i kön
Move down=Flytta ner
Move top=Flytta längst upp
Move up queue=Flytta till toppen av kön
Move up=Flytta upp
No updates have been found.~You are running the latest version of %s=Inga uppdateringar hittades.~Du kör senaste versionen av %s
Queue position=Köposition
Queue=Kö
Torrents that are idle for N minutes aren't counted toward the Download queue or Upload queue=Torrents som är inaktiva under N minuter räknas inte mot Download kön eller Upload kön
Tracker grouping=Trackergruppering
Upload queue size=Storlek på uppladdningskön
View=Visa
Visit home page=Besök hemsidan
days=dagar

Active time=Aktiv tid
Automatically add torrent links from the clipboard=Lägg automatiskt till torrent-länkar från urklipp
Copy file path to clipboard=Kopiera sökvägen till urklipp
Cumulative=Kumulativ
Current=Aktuell
Files added=Filer tillagda
Filter pane=Filterpanel
Global statistics=Global statistik
Info pane=Informationspanel
Statistics=Statistik
Status bar=Statusrad
%dd=%dd
%dh=%dh
%dm=%dm
All torrents=Alla torrents
Application options=Programalternativ
Ask for password=Fråga efter lösenord
Authentication required=Autentisering krävs
Average out transfer speeds to eliminate fluctuations=Jämna ut överföringshastigheten för att ta bort fluktuationer
Connect to %s=Anslut till %s
Connect to Transmission using proxy server=Anslut till Transmission via en proxyserver
Connect to Transmission=Anslut till Transmission
Connection name=Namn på anslutningen
Could not connect to tracker==Kunde inte ansluta till tracker
Data display=Datavisning
Data refresh interval when minimized=Uppdateringsintervall av data vid minimerad
Data refresh interval=Uppdateringsintervall av data
Default download folder on remote host=Nedladdningskatalog på Transmission-servern
Disconnect from Transmission=Stäng anslutningen till Transmission
Downloading torrent file=Laddar ner torrentfil
Font size=Storlek på typsnittet
Handle .torrent files by %s=Hantera .torrent-filer via %s
Handle magnet links by %s=Hantera magnetlänkar via %s
Invalid name specified=Felaktigt namn angivet
Manage connections to Transmission=Hantera anslutningar till Transmission
Manage connections=Hantera anslutningar
Network (WAN)=Nätverk (WAN)
New connection to Transmission=Ny anslutning till Transmission
Pick random port on Transmission launch=Använd slumpad port när Transmission startar
Please enter a password to connect to %s=Ange ett lösenord för att ansluta till %s
Please specify how %s will connect to a remote host running Transmission daemon (service)=Ange hur %s kommer ansluta till maskinen som kör Transmission-servern (service)
Prompt for download options when adding a new torrent=Fråga om nedladdningsalternativ när en ny torrent läggs till
RPC path=RPC-sökväg
Save as=Spara som
Seeding time=Uppladdningstid
Show advanced options=Visa avancerade alternativ
Show notifications in tray icon=Visa notifieringar i ikonen i aktivitetsfältet
System integration=Systemintegration
Torrent already exists in the list=Torrenten finns redan i listan
Torrent not registered with this tracker==Torrenten är inte registrerad hos denna tracker
Unable to find path mapping.~Use the application's options to setup path mappings=Hittar inte katalogen.~Använd inställningarna under alternativ för detta programmet för att justera katalogen (path)
Update trackers for the existing torrent?=Uppdatera trackers för den existerande torrenten?
You need to restart the application to apply changes=Du måste starta om programmet för att verkställa ändringarna
Development site=Webbplats för utveckling
Magnet Link=Magnetlänk
Status bar - Sizes=Statusrad - Storlekar
Total: %s=Totalt: %s
Remaining: %s=Kvarvarande: %s
Done: %s=Klart: %s
Selected: %s=Valt: %s
Export settings=Exportera inställningar
Import settings=Importera inställningar
Size left=Storlek kvar
Always auto-reconnect=Återanslut alltid automatiskt
The maximum history of directories for storage of torrents=Maximal historik över mappar för torrentlagring
Delete destination folder=Ta bort destinationsmapp
Template:=Mall:
for example: *.avi *.mkv tom*jerry*.avi=till exempel: *.avi *.mkv tom*jerry*.avi
Copy Magnet Link(s)=Kopiera magnetlänk(ar)
Application Options (Ctrl+F9)=Applikationsinställningar (Ctrl+F9)
Connection refused=Anslutning avvisad
Access violation=Åtkomstfel
Menu=Meny
Toolbar=Verktygsfält
Connection timed out=Anslutningstidsavbrott
Other Winsock error=Annat Winsock-fel
Default=Standard
Left->Right=Vänster->Höger
Right->Left=Höger->Vänster
Right->Left (No Align)=Höger->Vänster (ingen centrering)
Right->Left (Reading Only)=Höger->Vänster (endast läsning)
Host not found=Värden kunde inte hittas
User Menu=Användarmeny
Unauthorized User=Obehörig användare
