TranslationLanguage=Svenska

"Remote to local path mappings.~~Examples:~/share=\\pch\share~/var/downloads/music=Z:\music"="Mappning remote til lokala sökvägar.~~Till exempel:~/share=\\pch\share~/var/downloads/musik=Z:\musik"
%d x %s (have %d)=%d x %s (har %d)
%dd, %dh=%dd, %dh
%dh, %dm=%dh, %dm
%dm, %ds=%dm, %ds
%ds=%ds
%s (%d hashfails)=%s (%d checksummefel)
%s (%s done)=%s (%s klar)
'%s' has finished downloading='%s' är klar med nedladdningen
%s%s%d downloading, %d seeding%s%s, %s=%s%s%d laddar ned, %d delar%s%s, %s
&All=&Alla
&Close=&Stäng
&Help=&Hjälp
&Ignore=&Ignorera
&No=&Nej
&OK=&OK
&Open=&Öppna
&Retry=&Försök igen
&Save=&Spara
&Unlock=Lås upp
&Yes=&Ja
/s=/s
Abort=Avbryt
About=Om
Active=Aktiv
Add new torrent=Addera ny torrent
&Add torrent=Addera torrent
Added on=Adderades till
All=Alla
Are you sure to remove torrent '%s' and all associated DATA?=Är du säker på att du vill ta bort '%s' och alla tillhörande data?
Are you sure to remove torrent '%s'?=Är du säker på att du vill ta bort torrenten '%s'?
Authentication=Autentisering
b=b
Cancel=Avbryt
Client=Klient
Close to tray=Stäng till aktivitetsfältet
Comment=Kommentar
Completed on=Avslutad
Completed=Avslutad
Confirmation=Bekräftelse
Connect to daemon=Anslut till server
connected=Ansluten
Connecting to daemon=Ansluter till server
Connection error occurred=Anslutningsfel
Connection=Anslutning
Copy=Kopiera
Country=Land
Created on=Skapad
D: %s/s=D: %s/s
Delete host settings=Radera server inställningar
Destination folder=Destinationsmapp
Disconnected=Frånkopplad
Donate to support further development=Donera för att stödja fortsatt utveckling
Donate via PayPal,WebMoney,Credit card=Donera via PayPal,WebMoney,Credit card
Done=Färdig
Don't download=Ladda inte ned
Down limit=Ner gräns
Down speed=Nedladdningshastighet
Down=Ner
Download complete=Nedladdning klar
Download dir=Nedladdningsmapp
Download speed=Nedladdingshastighet
Downloaded=Nerladdad
Downloading=Laddar ner
Enable DHT=Aktivera DHT
Enable Peer Exchange=Aktivera Peer Exchange
Enable port forwarding=Aktivera portvidaresänding
Encryption disabled=Kryptering avstängd
Encryption enabled=Kryptering aktiverad
Encryption required=Kryptering krävs
Encryption=Kryptering
Error=Fel
ETA=ETA
E&xit=Avsluta
File name=Filnamn
Files=Filer
Finished=Avslutad
Flag images archive is needed to display country flags.~Download this archive now?=Ett arkiv med flaggbilder är nödvändigt för att visa landsflaggor.~Önskar du att ladda ned denna nu?
Flags=Flaggor
GB=GB
General=Allmänt
Geo IP database is needed to resolve country by IP address.~Download this database now?=En geo-IP databas är nödvändig för att visa vilket land en IP-adress tillhör.~Önskar du att ladda ned denna databasen nu??
Global bandwidth settings=Global bredbands inställningar
Global peer limit=Max antal globala kamrater
Hash=Checksum
Have=Ha
Hide=Dölj
High priority=Hög prioritet
high=hög
Host=värd
in swarm=i svärm
Inactive=Inaktiv
Incoming port is closed. Check your firewall settings=Inkommande port är stängd. Kontrollera brandväggs inställningarna
Incoming port tested successfully=Inkommande port är öppen
Incoming port=Inkommande port
Information=Information
Interface=Gränssnitt
KB/s=KB/s
KB=KB
Language=Språk
Last active=Senast aktiv
License=Licens
Low priority=Låg prioritet
low=låg
Max peers=Max antal peers
Maximum download speed=Max nedladdningshastighet
Maximum upload speed=Max uppladdningshastighet
MB=MB
Minimize to tray=Minimera till aktivitetsfältet
Name=Namn
No host name specified=Inget värdnamn specifierat
No proxy server specified=Ingen proxyserver specifierad
No to all=Nej till alla
Normal priority=Normal prioritet
normal=normal
of=av
OK=OK
Open containing folder=Öppna målmapp
Open=Öppna
Options=Alternativ
Password=Lösenord
Paths=Sökvägar
Pick random port on daemon launch=Välj en random port vid uppstart
Peer limit=Peer begränsning
Peers=Peers
Pieces=Delar
Port=Port
Priority=Prioritet
Properties=Egenskaper
Proxy password=Lösenord Proxy
Proxy port=Proxy port
Proxy server=Proxy server
Proxy user name=Användarnamn på proxy server
Ratio=Förhållande
Reconnect in %d seconds=Anslut på nytt om %d sekunder
Refresh interval=Uppdaterings intervall
Remaining=Återstående
Remote host=Fjärrserver
Remove torrent and Data=Ta bort torrent och data
Remove torrent=Ta bort torrent
Remove=Ta bort
Resolve country=Check land
Resolve host name=Check värdnamn
seconds=sekunder
Seed ratio=Delningsförhållande
Seeding=Delar
Seeds=Delare
Select a .torrent to open=Välj en .torrent att öppna
Select all=Välj alla
Select none=Välj ingen
Setup columns=Ställ in kolumner
Share ratio=Delningsförhållande
Show country flag=Visa flagga
Show parameters window when adding a new torrent=Visa parameterfönster när du lägger till en ny torrent
Show=Visa
Size=Storlek
skip=hoppa över
Start all torrents=Starta alla torrenter
Start torrent=Starta torrent
Start=Starta
Status=Status
Stop all torrents=Stoppa alla torrenter
Stop all=Stoppa alla
Stop torrent=Stopp torrent
Stop=Stopp
Stopped=Stoppad
TB=TB
Test port=Testa port
T&ools=Verktyg
Torrent contents=Innehåll i torrent
Torrent properties=Egenskaper för torrent
Torrent verification may take a long time.~Are you sure to start verification of torrent '%s'?=Torrentverifikation kan ta lång tid.~Är du säker på att du vill starta torrentverifikation '%s'?
&Torrent=Torrent
Torrents (*.torrent)|*.torrent|All files (*.*)|*.*=Torrenter (*.torrent)|*.torrent|Alla filar (*.*)|*.*
Total size=Total storlek
Tracker status=Trackerstatus
Tracker update on=Uppdaterar tracker
Tracker=Tracker
Trackers=Trackers
Transfer=Överföring
Transmission options=Alternativ för Transmission
Transmission%s at %s:%s=Transmission%s på %s:%s
Tray icon always visible=Ikon i aktivitetsfältet alltid synlig
Tray icon=Ikon i aktivitetsfältet
U: %s/s=U: %s/s
Unable to extract flag image=Kunde inte hämta flaggbild
Unable to find path mapping.~Use program's options to setup path mappings=Kunde inte finna servermappen lokalt.~Använd programmets alternativ för att ställa in server till klientens mapprelationer
Unable to get files list=Kunde inte finna fillista
Unknown=Okänt
Up limit=Uppladdnings gräns
Up speed=Uppladdnings hastighet
Up=Upp
Update complete=Uppdatering genomförd
Update GeoIP database=Uppdatera GeoIP databas
Update in=Uppdaterar om
Updating=Uppdaterar
Upload speed=Uppladdnings hastighet
Uploaded=Uppladdat
Use proxy server=Använd proxyserver
User name=Användarnamn
Verify torrent=Verifiera torrents
&Verify=Verifiera
Verifying=Verifierar
Version %s=Version %s
Waiting=Väntar
Warning=Varning
Wasted=Bortkastad
Working=Arbetar
Yes to &All=Ja till &Alla
You should restart the application to apply changes=Du måste starta om programmet för att ändringarna ska träda i kraft
No tracker=Ingen tracker
Tracker did not respond=Trackern svarade inte
%s downloaded=%s nedladdat
%s of %s downloaded=%s av %s nedladdad
%d torrents=%d torrents
Add .part extension to incomplete files=Lägg till .part på ofullständiga filer
Add torrent link=Lägg till en torrentlänk
Are you sure to remove %d selected torrents and all their associated DATA?=är du säker på att du önskar att ta bort %d valda torrenter och alla tilhörande data?
Are you sure to remove %d selected torrents?=är du säker på att du önskar att ta bort %d valda torrenter?
Bandwidth=Bandbredd
Directory for incomplete files=Mapp för ofullständiga filer
Download=Ladda ner
Enable blocklist=Aktivera blockeringslistan
ID=ID
Move torrent data from current location to new location=Flytta data från nuvarande till ny plats
Network=Nätverk
New location for torrent data=Ny plats för torrent data
No link was specified=Ingen länk specifierad 
No torrent location was specified=Ingen torrentplats var specifierad
Path=Sökväg
Reannounce (get more peers)=Tillkännage (skaffa flera peers)
Set data location=Sätt dataplats
Size to download=Storlek på nedladdning
The block list has been updated successfully.~The list entries count: %d=Blockeringslistan blev uppdaterad.~Det är %d registrerade i listan
The directory for incomplete files was not specified=Mappen för ofullständiga filer var inte specifierad
The downloads directory was not specified=Det blev inte specifierat en neddladdnings map
Torrent data location=Dataplats for torrent
Torrents=Torrents
Unable to execute "%s"=Kunde inte köra "%s"
Update blocklist=Uppdatera blockeringslista
URL of a .torrent file or a magnet link=Adressen till en .torrent-fil eller en magnet-länk
Columns setup=Kolumn inställning
Add torrent=Lägg till torrent
Delete a .torrent file after after a successful addition=Ta bort .torrent-filen efter att den är uppladdad till servern
Torrent=Torrent
Torrents verification may take a long time.~Are you sure to start verification of %d torrents?=Dataverifiering kan ta lång tid.~Är du säker på att du önskar att verifiera %d torrenter?
Unable to load OpenSSL library files: %s and %s=Klarade inte att ladda OpenSSL biblioteks filerna: %s och %s från OpenSSL
Use SSL=Använd SSL
Add tracker=Lägg till tracker
Alternate bandwidth settings=Alternativ bandbredds inställingar
Apply alternate bandwidth settings automatically=Använd alternativ bandbreds inställningar automatiskt
Are you sure to delete connection '%s'?=Är du säker på att du vill ta bort anslutningen '%s'?
Are you sure to remove tracker '%s'?=Är du säker på att du vill ta bort trackern '%s'?
Connection options=Anslutnings inställningar
Days=Dagar
Delete=Ta bort
Disconnect=Koppla från
Disk cache size=Storlek på disk cachen
Download speeds (KB/s)=Nedladdingshastighet (KB/s)
Edit tracker=Redigera tracker
Enable Local Peer Discovery=Aktivera Lokal Peer upptäckt
Free disk space=Ledigt diskutrymme
Free: %s=Ledigt: %s
From=Från
minutes=minuter
Misc=Diverse
New connection=Ny anslutning
New=Ny
No tracker URL was specified=Ingen Trackeradress var specifierad
Proxy=Proxy
Refresh interval when minimized=uppdateringsfrekvens vid minimerad
Remove tracker=Radera tracker
Rename=Byt namn
Speed limit menu items=Hastighetsbegränsningar
Stop seeding when inactive for=Avsluta delning när inaktiv i
The blocklist URL was not specified=Adressen till blockeringslistan ej angiven
The invalid time value was entered=Ett ogiltig tidsvärde angavs
to=till
Tracker announce URL=Trackerns annonseringsadress
Tracker properties=Trackerinställningar
Unlimited=Obegränsat
Upload speeds (KB/s)=Uppladdnings hastighet (KB/s)
Use alternate bandwidth settings=Använd alternativ bandbredds inställning
average=genomsnitt
Browse=Bläddra
Enable µTP=Aktivera µTP
Select a folder for download=Välj nedladdningsmapp
Select torrent location=Välj torrentplats
A new version of %s is available.~Your current version: %s~The new version: %s~~Do you wish to open the Downloads web page?=A new version of %s is available.~Your current version: %s~The new version: %s~~Do you wish to open the Downloads web page?
Advanced=Avancerad
Check for new version every=Sök efter nya versioner varje
Check for updates=Sök efter uppdateringar
Consider active torrents as stalled when idle for=Consider active torrents as stalled when idle for
Do you wish to enable automatic checking for a new version of %s?=Vill du aktivera automatisk kontroll av nya versioner av %s?
Donate!=Donera!
Download queue size=Storlek på download kön
Error checking for new version=Fel kontroll av ny version
Folder grouping=Gruppering av mappar
Force start=Tvinga start
Home page=Hemsida
Modify trackers=Modifiera trackers
Move bottom=Flytta till botten av kön
Move down queue=Flytta ner i kön
Move down=Flytta ner
Move top=Flytta längst upp
Move up queue=Flytta till toppen av kön
Move up=Flytta upp
No updates have been found.~You are running the latest version of %s=Inga uppdateringar hittades.~Du kör senaste versionen av %s
Queue position=Kö position
Queue=Kö
Torrents that are idle for N minuets aren't counted toward the Download queue or Upload queue=Torrents som är inaktiva under N minuter räknas inte mot Download kön eller Upload kön
Tracker grouping=Tracker gruppering
Upload queue size=Upload kö storlek
User interface scaling=Användargränssnitt skalning
View=Visa
Visit home page=Besök hemsidan
days=dagar

Active time=Active time
Automatically add torrent links from the clipboard=Automatically add torrent links from the clipboard
Copy file path to clipboard=Copy file path to clipboard
Cumulative=Cumulative
Current=Current
Files added=Files added
Filter pane=Filter pane
Global statistics=Global statistics
Info pane=Info pane
Statistics=Statistics
Status bar=Status bar
